module forwarding_logic (IFETCH_instruction, REG_instruction, EXEC_instruction);
	input logic [31:0] IFETCH_instruction, REG_instruction, EXEC_instruction;
	always_comb begin
		
	end

endmodule 