module Execute (op_result, mem_wr, reg_wr, mem_to_reg, Rd);

endmodule 