module RegisterFetch (Da, Db, Rd, mem_wr, reg_wr, alu_src, ctrl, mem_to_reg, setFlags, shift, imm_or_D9, D9, Imm12,
							 REG_Da, REG_Db, REG_Rd, REG_mem_wr, REG_reg_wr, REG_alu_src, REG_ctrl, REG_mem_to_reg, REG_setFlags, REG_shift, REG_imm_or_D9, REG_D9, REG_Imm12);
	// finish later

endmodule 